package pkg_alu;
  typedef enum logic [3:0] {
  	A_ADD ,
  	A_SUB ,
  	A_SLT ,
  	A_SLTU,
  	A_XOR ,
  	A_OR  ,
  	A_AND ,
  	A_SLL ,
  	A_SRL ,
  	A_SRA ,
  	A_LUI
  } alu_op_e;

endpackage

